`timescale 1ns / 1ps
`default_nettype none
`default_nettype wire



module controller (
    input wire [2:0] opcode,
    
)

endmodule