`define BUS_WIDTH 7



// A register file meant to supply values to a tensor core.
// This register file exposes all of the wires to each register, so a tensor core can take each of the values inside the registers in a single clock cycle 
module tensor_core_register_file (
    input logic clock_in,
    input logic reset_in,

    // writing elements 4 at a time
    input logic quad_write_enable_in,
    input logic [2:0] quad_write_register_address_in, // supports values 0 to 4
    input logic signed [`BUS_WIDTH:0] quad_write_data_in [4],

    // bulk read
    output logic signed [`BUS_WIDTH:0] bulk_read_data_out [2] [3] [3]
);


    reg signed [7:0] registers [2] [3] [3];



    always_comb begin

        // assign bulk read wires
        for (int n = 0; n < 2; n++) begin
            for (int i = 0; i < 3; i++) begin
                for (int j = 0; j < 3; j++) begin
                    bulk_read_data_out[n][i][j] = registers[n][i][j];
                end
            end
        end

    end


    always_ff @(posedge clock_in) begin

        // quad write
        if (quad_write_enable_in && reset_in == 0) begin
            for (int i = 0; i < 4; i++) begin
                registers[((quad_write_register_address_in<<2)+i)/9][(((quad_write_register_address_in<<2)+i)%9)/3][((quad_write_register_address_in<<2)+i)%3] <= quad_write_data_in[i];
            end
        end

        // reset logic
        else if (reset_in == 1) begin
            for (int i = 0; i < 2; i++) begin
                for (int j = 0; j < 3; j++) begin
                    for (int k = 0; k < 3; k++) begin
                        registers[i][j][k] <= 0;
                    end
                end
            end
        end
    end



    // // make the registers visible to gtkwave
    // genvar i, j, k;
    // generate
    //     for (i = 0; i < 2; i++) begin : expose_regs1
    //         for (j = 0; j < 3; j++) begin : expose_regs2
    //             for (k = 0; k < 3; k++) begin : expose_regs3
    //                 wire [`BUS_WIDTH:0] reg_wire = registers[i][j][k];
    //                 wire [`BUS_WIDTH:0] bulk_read_data_out_ = bulk_read_data_out[i][j][k];
    //                 wire [`BUS_WIDTH:0] bulk_write_data_in_ = bulk_write_data_in[i][j][k];
    //             end
    //         end
    //     end
    // endgenerate


endmodule