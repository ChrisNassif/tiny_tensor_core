`timescale 1ns / 1ps
`default_nettype none
`default_nettype wire


module program_counter(
    output [7:0] program_counter_out;
)

endmodule